module sort